netcdf s117e {
// Program to define the netcdf structure of Phil Morgan's example
// which uses the data in s117e.mat.

dimensions:
   depths = 32, lat = 127, lon = 127;

variables:
   float gvel(depths,lat);
      gvel:long_name       = "geostrophic velocity";
      gvel:units           = "m/sec";
      gvel:_FillValue      = -9.99e+2f;
      gvel:missing_value   = -9.99e+2f;

   float sal(depths,lat);
      sal:long_name       = "salinity";
      sal:units           = "ppt";
      sal:_FillValue      = -9.99e+2f;
      sal:missing_value   = -9.99e+2f;

   float theta(depths,lat);
      theta:long_name       = "potential temperature";
      theta:units           = "degrees celsius";
      theta:_FillValue      = -9.99e+2f;
      theta:missing_value   = -9.99e+2f;

   float depths(depths);
      depths:long_name       = "depth for sample";
      depths:units           = "meters";


   float lat(lat);
      lat:long_name       = "latitude for sample";
      lat:units           = "degrees north";


   float lon(lon);
      lon:long_name       = "longitude for sample";
      lon:units           = "degrees east";

// global attributes

:source = "Phil Morgan - example file in s117e.mat";
:title = "Oceanographic data from a 117E meridional section";
:history = "netCDF file created by Jim Mansbridge";
}